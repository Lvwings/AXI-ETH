         
//----------AXIS PARAMETERS-------------------

                  
            
// IP datagram header format
//
//      0          4          8                      16      19             24                    31
//      --------------------------------------------------------------------------------------------
//      | Version  | *Header  |    Service Type      |        Total Length including header        |
//      |   (4)    |  Length  |     (ignored)        |                 (in bytes)                  |
//       ///////////*IP_VS_LEN_TOS*//////////////////////////////// *TX_IP_TOTAL_LEN*///////////////
//      --------------------------------------------------------------------------------------------
//      |           Identification                   | Flags |       Fragment Offset               |
//      |                                            |       |      (in 32 bit words)              |
//      //////////////*IP_IDENTIF*////////////////////////////////*IP_FLAG_OFFSET*//////////////////
//      --------------------------------------------------------------------------------------------
//      |    Time To Live     |       Protocol       |             Header Checksum                 |
//      |     (ignored)       |                      |                                             |
//      ////////////////*IP_TTL_PROTO*//////////////////////////////*TX_IP_HEADER_CKS*//////////////
//      --------------------------------------------------------------------------------------------
//      |                                   Source IP Address                                      |
//      |                                ////////*IP_SA*/////////                                  |
//      --------------------------------------------------------------------------------------------
//      |                                 Destination IP Address                                   |
//      |                                ////////*IP_DA*/////////                                  |
//      --------------------------------------------------------------------------------------------
//      |                          Options (if any - ignored)               |       Padding        |
//      |                                                                   |      (if needed)     |
//      --------------------------------------------------------------------------------------------
//      |                                          Data                                            |
//      |                                                                                          |
//      --------------------------------------------------------------------------------------------
//      |                                          ....                                            |
//      |                                                                                          |
//      --------------------------------------------------------------------------------------------
//
// * - in 32 bit words
           
localparam  PREAMBLE_REG   =   64'h5555_5555_5555_55d5,    //  前导码
            PREAMBLE_WORD  =   8'd8,
            //------------以太网首部-----------------       //  000a_3501_fec0_ffff_ffff_ffff_0800
            IP_TYPE        =   16'h0800,                   //  IP帧
            ARP_TYPE       =     16'h0806,                           //    ARP帧
            ETH_WORD       =   8'd14,
            //-------------IP首部----------------------     //  4500_0014_0000_4000_8011_c0a8_0003_c0a8_0002
            IP_VS_LEN_TOS  =   16'h4500,                   //  IP版本(4)+首部长度(20)+服务类型
            IP_FLAG_OFFSET =   16'h4000,                   //  IP标志+帧偏移
            IP_TTL         =   8'h80,                      //  IP帧生存时间
            UDP_PROTO      =   8'h11,                                // UDP协议
            ICMP_PROTO     =     8'h01,                                    // ICMP协议
            IP_WORD        =   8'd20,
            //-------------UDP首部---------------------     //  1F90_1F90_0010_3F30
            UDP_WORD       =   8'd8, 
            //-------------等待---------------------
            WAIT_DEADLINE  =     9'd100,
            //-------------数据---------------------
            FLAG_MOTOR     =     32'hE1EC_0C0D,
            FLAG_AD        =     32'hAD86_86DA,
            FLAG_WORD      =     8'd4,
            MOTOR_WORD     =     8'd38,
            AD_WORD        =     8'd128,
            //-------------ARP---------------------
            ARP_HEAD       =     64'h0001_0800_0604_0002,      //硬件类型+协议类型+硬件地址长度+协议地址长度+操作字段
            ARP_WORD       =     8'd48,                                    // 28 + 20 ->有20位填充数据FF
            ARP_REQUEST    =     16'h0001,
            //-------------ICMP---------------------
            PING_REQ       =     8'h08,
            ICMP_TYPE      =     8'h00,
            ICMP_CODE      =     8'h00,
            ICMP_WORD      =     8'd40,                  
            //-------------CRC---------------------
            CRC_WORD       =   8'd4;
//---------------------------------------
