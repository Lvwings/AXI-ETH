// IP datagram header format
//
//      0          4          8                      16      19             24                    31
//      --------------------------------------------------------------------------------------------
//      | Version  | *Header  |    Service Type      |        Total Length including header        |
//      |   (4)    |  Length  |     (ignored)        |                 (in bytes)                  |
//      --------------------------------------------------------------------------------------------
//      |           Identification                   | Flags |       Fragment Offset               |
//      |                                            |       |      (in 32 bit words)              |
//      --------------------------------------------------------------------------------------------
//      |    Time To Live     |       Protocol       |             Header Checksum                 |
//      |     (ignored)       |                      |                                             |
//      --------------------------------------------------------------------------------------------
//      |                                   Source IP Address                                      |
//      |                                                                                          |
//      --------------------------------------------------------------------------------------------
//      |                                 Destination IP Address                                   |
//      |                                                                                          |
//      --------------------------------------------------------------------------------------------
//      |                          Options (if any - ignored)               |       Padding        |
//      |                                                                   |      (if needed)     |
//      --------------------------------------------------------------------------------------------
//      |                                          Data                                            |
//      |                                                                                          |
//      --------------------------------------------------------------------------------------------
//      |                                          ....                                            |
//      |                                                                                          |
//      --------------------------------------------------------------------------------------------
//
// * - in 32 bit words

localparam  PREAMBLE_REG  =   64'h5555_5555_5555_55d5,    //  前导码
            PREAMBLE_WORD =   8'd8,
            //------------以太网首部-----------------       //  000a_3501_fec0_ffff_ffff_ffff_0800
            IP_TYPE       =   16'h0800,                   //  IP帧
            ARP_TYPE      =   16'h0806,                           //    ARP帧
            ETH_WORD      =   8'd14,
            //-------------IP首部----------------------     //  4500_0014_0000_4000_8011_c0a8_0003_c0a8_0002
            UDP_PROTO     =   8'h11,                                // UDP协议
            ICMP_PROTO    =   8'h01,                                    // ICMP协议
            IP_WORD       =   8'd20,
            //-------------UDP首部---------------------     //  1F90_1F90_0010_3F30
            UDP_WORD      =   8'd8,                       
            //-------------数据---------------------
            FLAG_MOTOR    =   32'hE1EC_0C0D,              //   电机配置固定标识
            DATA_WORD     =   8'd44,                                  // 30字节数据 + 最后两位填充
            //-------------ARP---------------------
            ARP_WORD      =   8'd28,                  //    28 + 18 18 位00填充
            ARP_REQUEST   =   16'h0001,
            //-------------ICMP---------------------
            PING_REQ      =   8'h08,
            ICMP_WORD     =   8'd40,
            //-------------CRC---------------------
            CRC_WORD      =   8'd4;